module cpu_tb;

    parameter TIMEOUT_CYCLES = 10000;

    logic clk;
    logic reset;

    logic active;
    logic [31:0] register_v0;

    logic clk_enable;

    logic[3:0] instr_address;
    logic[31:0] instr_readdata;


    logic[3:0]  data_address;
    logic        data_write;
    logic        data_read;
    logic[31:0]  data_writedata;
    logic[31:0]  data_readdata;

    RAM_32x4GB ramInst(clk, instr_address, instr_readdata);

    RAM_32x8_delay0 ramDataInst(clk, data_address, data_write, data_read, data_writedata, data_readdata);
    
    mips_cpu_harvard cpuInst(clk, reset, active, register_v0, clk_enable, instr_address, instr_readdata, data_address, data_write, data_read, data_writedata, data_readdata);

    // Generate clock
    initial begin
        $dumpfile("cpu.vcd");
        $dumpvars(0, cpu_tb);
        clk=0;
        //data_readdata=32'b00000000000000000000000111111101;
        repeat (TIMEOUT_CYCLES) begin
            #10;
            clk = !clk;
            #10;
            clk = !clk;
        end

        $fatal(2, "Simulation did not finish within %d cycles.", TIMEOUT_CYCLES);
    end

    initial begin
        reset <= 0;

        @(posedge clk);
        reset <= 1;

        @(posedge clk);
        reset <= 0;
        $display("reset back to 0");

        @(posedge clk);
        if(active==1) $display("active set to 1");
        else $display("TB : CPU did not set running=1 after reset.");


        while (active) begin
            @(posedge clk);
        end

        $display("TB : finished; running=0");
        $display("register_v0 value: %d ", register_v0);
        $finish;
        
    end

    

endmodule